# ====================================================================
#
#      can_loop.cdl
#
#      eCos CAN LOOP configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Uwe Kindler
# Original data:  gthomas
# Contributors:
# Date:           2005-07-11
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_CAN_LOOP {
    display       "Loop CAN device drivers"

    parent        CYGPKG_IO_CAN_DEVICES
    active_if     CYGPKG_IO_CAN
    requires      CYGPKG_ERROR
    include_dir   cyg/io
    include_files ; # none _exported_ whatsoever

    description   "
       This package contains the loop CAN device driver."

    compile       -library=libextras.a loop_can.c

    # Support up to two CAN loop device.
    for { set ::loopcan 0 } { $::loopcan < 2 } { incr ::loopcan } {
    
    cdl_component CYGPKG_DEVS_CAN_LOOP_CAN[set ::loopcan] {
        display       "LOOP CAN channel [set ::loopcan] driver"
        flavor        bool
        default_value 0
        implements    CYGINT_IO_CAN_TIMESTAMP
        implements    CYGINT_IO_CAN_TX_EVENTS
        implements    CYGINT_IO_CAN_STD_CAN_ID
        implements    CYGINT_IO_CAN_EXT_CAN_ID
        description   "
            This option includes the CAN loop device driver for channel [set ::loopcan]." 
    
        cdl_option CYGDAT_DEVS_CAN_LOOP_CAN[set ::loopcan]_NAME {
            display       "Device name for LOOP CAN channel [set ::loopcan]"
            flavor        data
            default_value [format {"\"/dev/can%d\""} $::loopcan]
            description   "
                This option specifies the device name for loop CAN channel [set ::loopcan]."
        }
    
        cdl_option CYGNUM_DEVS_CAN_LOOP_CAN[set ::loopcan]_KBAUD {
            display       "Baud rate for the LOOP CAN channel [set ::loopcan] driver"
            flavor        data
            default_value   100
                legal_values    { 10 20 50 100 125 250 500 800 1000 }
                description "This option determines the initial baud rate in KBaud for 
                             loop CAN channel [set ::loopcan]."
        }
        
        cdl_option CYGNUM_DEVS_CAN_LOOP_CAN[set ::loopcan]_QUEUESIZE_TX {
                display     "Size of TX Queue for loop CAN channel [set ::loopcan]"
                flavor      data
                default_value   32
                legal_values    16 to 512
                description "
                    The CAN device driver will run in interrupt mode and will
                    perform buffering of outgoing data. This option controls the number
                    of CAN messages the TX queue can store."
            }
            
            cdl_option CYGNUM_DEVS_CAN_LOOP_CAN[set ::loopcan]_QUEUESIZE_RX {
                display     "Size of RX Queue for the loop CAN channel [set ::loopcan]"
                flavor      data
                default_value   32
                legal_values    16 to 512
                description "
                    The CAN device driver will run in interrupt mode and will
                    perform buffering of incoming data. This option controls the number
                    of CAN events the RX queue can store."
            }
        }
    }
    

    cdl_component CYGPKG_DEVS_CAN_LOOP_OPTIONS {
        display "CAN device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."

        
        cdl_option CYGPKG_DEVS_CAN_LOOP_TESTS {
            display "CAN loop device driver tests"
            flavor  data
            calculated { "tests/can_rdwr tests/can_timeout tests/can_txevent tests/can_overrun1 tests/can_overrun2 tests/can_nonblock tests/can_callback" }         
            description   "
                This option specifies the set of tests for the CAN loop device drivers."
        }
    }
}

# EOF can_loop.cdl
